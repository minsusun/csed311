module immediate_generator(
    input part_of_inst,
    output imm_gen_out
);

endmodule
