// Do not submit this file.
module top(input reset,
           input clk,
           output is_halted,
           output [31:0] print_reg [0:31]);

  cpu cpu(
    .reset(reset), 
    .clk(clk),
    .is_halted(is_halted),
    .print_reg(print_reg)
  );

endmodule
