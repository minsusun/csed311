module alu_control_unit(
    input part_of_inst,
    output alu_op
);

endmodule
